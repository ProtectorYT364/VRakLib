module protocol

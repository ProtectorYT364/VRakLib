module vraklib

import net
import time
import bstone

pub struct VRakLib {
pub mut:
	address              net.Addr
	session_manager      SessionManager
	shutdown             bool
	pong_data PongData
}

pub fn new_vraklib(shared config bstone.ServerConfig) &VRakLib {//TODO pass server config for pongdata
	address := rlock config{
		config.addr
	}
	pongdata := PongData{
		server_id: server_guid
		port: address.port
	}
	vr := &VRakLib{
		address: address
		pong_data: pongdata
	}
	return vr
}

pub fn (mut r VRakLib) start(shared logger bstone.Log) {
	println('RakLib thread starting on $r.address')
	socket := create_socket(r.address) or { panic(err) }

	mut session_manager := new_session_manager(r, socket)
	r.session_manager = session_manager
	session_manager.start(shared logger)//TODO check if this blocks
	session_manager.stop()
	println('Shutdown raklib? $r.shutdown')
	r.stop()
}

pub fn (mut r VRakLib) stop() {
	println('Shutting down RakLib')
	r.shutdown = true
	r.session_manager.stop()
}

// timestamp returns a timestamp in milliseconds.
pub fn timestamp() u64 {
	return time.now().unix_time_milli()
}
module vraklib

pub struct InternetAddress {
pub mut:
    ip string
    port u16
    version byte
}

module vraklib

module vraklib

pub type U24 = u32

pub fn u32(u U24) u32{
	return u
}

pub fn u24<T>(u T) U24{
	return u
}